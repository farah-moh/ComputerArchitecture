Library IEEE;
use IEEE.std_logic_1164.all;


entity tb_PartB is
end entity;


Architecture testingPartB of tb_PartB is

component PartB is 
port  (
    A :    in std_logic_vector(15 downto 0); 
    B:     in std_logic_vector(15 downto 0); 
    sel :     in std_logic_vector (1 downto 0);
    Cin:    in std_logic;
    Cout :     out std_logic;
    F :     out std_logic_vector(15 downto 0)
);
end component;

Signal test_A:      std_logic_vector(15 downto 0);
Signal test_B:      std_logic_vector(15 downto 0);
Signal test_sel:    std_logic_vector (1 downto 0);
Signal test_Cin:    std_logic;
Signal test_Cout:   std_logic;
Signal test_F:      std_logic_vector(15 downto 0);

Begin

  U1: PartB port map (test_A,test_B,test_sel,test_Cin,test_Cout,test_F);
process
begin

test_Cin    <= '0';

-- test case 1:
test_A      <= x"F000";
test_B      <= x"00B0";
test_sel    <= "00";

wait for 10 ns;

assert (test_F=x"F0B0")
    report "Failed Case: " & to_hstring(test_A) &" " & to_hstring(test_B) &" "& to_hstring(test_sel) &" "& std_logic'image(test_Cin) & " output: " & to_hstring(test_F)  severity error;

-- test case 2:
test_A      <= x"F000";
test_B      <= x"000B";
test_sel    <= "01";

wait for 10 ns;

assert (test_F=x"0000")
    report "Failed Case: " & to_hstring(test_A) &" " & to_hstring(test_B) &" "& to_hstring(test_sel) &" "& std_logic'image(test_Cin) & " output: " & to_hstring(test_F)  severity error;

-- test case 3:
test_A      <= x"F000";
test_B      <= x"B000";
test_sel    <= "10";

wait for 10 ns;

assert (test_F=x"0FFF")
    report "Failed Case: " & to_hstring(test_A) &" " & to_hstring(test_B) &" "& to_hstring(test_sel) &" "& std_logic'image(test_Cin) & " output: " & to_hstring(test_F)  severity error;

-- test case 4:
test_A      <= x"F000";
test_B      <= x"0000";
test_sel    <= "11";

wait for 10 ns;

assert (test_F=x"0FFF")
    report "Failed Case: " & to_hstring(test_A) &" " & to_hstring(test_B) &" "& to_hstring(test_sel) &" "& std_logic'image(test_Cin) & " output: " & to_hstring(test_F)  severity error;


wait for 10 ns;
report "Done";
wait;



end process;



end testingPartB;
